
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


USE IEEE.NUMERIC_STD.ALL;

ENTITY SEVSEG_DRIVER IS
    PORT ( D8: IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
           D7 : IN  STD_LOGIC_vector (3 DOWNTO 0);
			  D6 : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			  D5 : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			  D4 : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			  D3 : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			  D2 : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			  D1  : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
           CLK : IN  STD_LOGIC;
			  SEV_SEG_DATA : OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
           SEV_SEG_DRIVER : OUT  STD_LOGIC_VECTOR (7 DOWNTO 0)
			  );
END SEVSEG_DRIVER;

ARCHITECTURE BEHAVIORAL OF SEVSEG_DRIVER IS

SIGNAL COUNTER : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";

BEGIN

---mods

--INCREMENT COUNTER
PROCESS_CLK : PROCESS(CLK)
BEGIN
	IF(CLK'EVENT AND CLK = '1') THEN
			COUNTER <= COUNTER + 1;
			IF(COUNTER = "111" )THEN
			 COUNTER <= "000";
			END IF;
	END IF;
END PROCESS;

-- SEV_SEG DATA
WITH COUNTER SELECT SEV_SEG_DATA <=

	D8 WHEN "000",
	D7 WHEN "001",
	D6 WHEN "010",
	D5 WHEN "011",
	D4 WHEN "100",
	D3 WHEN "101",
	D2 WHEN "110",
	D1 WHEN "111",
	"1001" WHEN OTHERS; 
--DATA END

--SEV_SEG_CONTROLLER
WITH COUNTER SELECT SEV_SEG_DRIVER <=
"01111111" WHEN "000", 
"10111111" WHEN "001", 
"11011111" WHEN "010", 
"11101111" WHEN "011", 
"11110111" WHEN "100", 
"11111011" WHEN "101",
"11111101" WHEN "110",
"11111110" WHEN "111",
"00001111" WHEN OTHERS;
--SEV_SEG CONTROLLER END

END BEHAVIORAL;

