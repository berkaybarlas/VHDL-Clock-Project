
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY SEVSEG_DECODER IS
    PORT ( INPUT : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
           SEVSEG_BUS : OUT  STD_LOGIC_VECTOR (6 DOWNTO 0));
END SEVSEG_DECODER;

ARCHITECTURE BEHAVIORAL OF SEVSEG_DECODER IS

BEGIN

WITH INPUT SELECT SEVSEG_BUS <=
	"0000001" when "0000", --0
	"1001111" when "0001", --1
	"0010010" when "0010", --2
	"0000110" when "0011", --3
	"1001100" when "0100", --4
	"0100100" when "0101", --5
	"0100000" when "0110", --6
	"0001111" when "0111", --7
	"0000000" when "1000", --8
	"0000100" when "1001", --9
	
	"0001000" when "1010", --A
	"0110001" when "1011", --C
	"1100010" when "1100", --O
	"1110001" when "1101", --L
	"1111010" when "1111", --R
	"1001000" when "1110", --H
	
	

	"0000100" WHEN OTHERS;
END BEHAVIORAL;

